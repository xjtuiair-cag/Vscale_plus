`define N_EXT_INTS 8